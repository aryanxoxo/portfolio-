
`default_nettype none
module simple_ipod_solution(

    //////////// CLOCK //////////
    CLOCK_50,

    //////////// LED //////////
    LEDR,

    //////////// KEY //////////
    KEY,

    //////////// SW //////////
    SW,

    //////////// SEG7 //////////
    HEX0,
    HEX1,
    HEX2,
    HEX3,
    HEX4,
    HEX5,

    //////////// Audio //////////
    AUD_ADCDAT,
    AUD_ADCLRCK,
    AUD_BCLK,
    AUD_DACDAT,
    AUD_DACLRCK,
    AUD_XCK,

    //////////// I2C for Audio  //////////
    FPGA_I2C_SCLK,
    FPGA_I2C_SDAT,
    
    
    //////// PS2 //////////
    PS2_CLK,
    PS2_DAT,
    
    //////// SDRAM //////////
    DRAM_ADDR,
    DRAM_BA,
    DRAM_CAS_N,
    DRAM_CKE,
    DRAM_CLK,
    DRAM_CS_N,
    DRAM_DQ,
    DRAM_LDQM,
    DRAM_UDQM,
    DRAM_RAS_N,
    DRAM_WE_N,
    
    //////// GPIO //////////
    GPIO_0,
    GPIO_1
    
);
`define zero_pad(width,signal)  {{((width)-$size(signal)){1'b0}},(signal)}
//=======================================================
//  PORT declarations
//=======================================================

//////////// CLOCK //////////
input                       CLOCK_50;

//////////// LED //////////
output           [9:0]      LEDR;

//////////// KEY //////////
input            [3:0]      KEY;

//////////// SW //////////
input            [9:0]      SW;

//////////// SEG7 //////////
output           [6:0]      HEX0;
output           [6:0]      HEX1;
output           [6:0]      HEX2;
output           [6:0]      HEX3;
output           [6:0]      HEX4;
output           [6:0]      HEX5;



//////////// Audio //////////
input                       AUD_ADCDAT;
inout                       AUD_ADCLRCK;
inout                       AUD_BCLK;
output                      AUD_DACDAT;
inout                       AUD_DACLRCK;
output                      AUD_XCK;

//////////// I2C for Audio  //////////
output                      FPGA_I2C_SCLK;
inout                       FPGA_I2C_SDAT;

//////////// PS2 //////////
inout                       PS2_CLK;
inout                       PS2_DAT;

//////////// GPIO //////////
inout           [35:0]      GPIO_0;
inout           [35:0]      GPIO_1;
                
                
//////////// SDRAM //////////
output          [12:0]      DRAM_ADDR;
output        [1:0]         DRAM_BA;
output                      DRAM_CAS_N;
output                      DRAM_CKE;
output                      DRAM_CLK;
output                      DRAM_CS_N;
inout           [15:0]      DRAM_DQ;
output                      DRAM_LDQM;
output                      DRAM_UDQM;
output                      DRAM_RAS_N;
output                      DRAM_WE_N;


//=======================================================
//  REG/WIRE declarations
//=======================================================
// Input and output declarations
logic CLK_50M;
logic  [7:0] LED;
assign CLK_50M =  CLOCK_50;
assign LEDR[7:0] = LED[7:0];

//Character definitions

//numbers
parameter character_0 =8'h30;
parameter character_1 =8'h31;
parameter character_2 =8'h32;
parameter character_3 =8'h33;
parameter character_4 =8'h34;
parameter character_5 =8'h35;
parameter character_6 =8'h36;
parameter character_7 =8'h37;
parameter character_8 =8'h38;
parameter character_9 =8'h39;


//Uppercase Letters
parameter character_A =8'h41;
parameter character_B =8'h42;
parameter character_C =8'h43;
parameter character_D =8'h44;
parameter character_E =8'h45;
parameter character_F =8'h46;
parameter character_G =8'h47;
parameter character_H =8'h48;
parameter character_I =8'h49;
parameter character_J =8'h4A;
parameter character_K =8'h4B;
parameter character_L =8'h4C;
parameter character_M =8'h4D;
parameter character_N =8'h4E;
parameter character_O =8'h4F;
parameter character_P =8'h50;
parameter character_Q =8'h51;
parameter character_R =8'h52;
parameter character_S =8'h53;
parameter character_T =8'h54;
parameter character_U =8'h55;
parameter character_V =8'h56;
parameter character_W =8'h57;
parameter character_X =8'h58;
parameter character_Y =8'h59;
parameter character_Z =8'h5A;

//Lowercase Letters
parameter character_lowercase_a= 8'h61;
parameter character_lowercase_b= 8'h62;
parameter character_lowercase_c= 8'h63;
parameter character_lowercase_d= 8'h64;
parameter character_lowercase_e= 8'h65;
parameter character_lowercase_f= 8'h66;
parameter character_lowercase_g= 8'h67;
parameter character_lowercase_h= 8'h68;
parameter character_lowercase_i= 8'h69;
parameter character_lowercase_j= 8'h6A;
parameter character_lowercase_k= 8'h6B;
parameter character_lowercase_l= 8'h6C;
parameter character_lowercase_m= 8'h6D;
parameter character_lowercase_n= 8'h6E;
parameter character_lowercase_o= 8'h6F;
parameter character_lowercase_p= 8'h70;
parameter character_lowercase_q= 8'h71;
parameter character_lowercase_r= 8'h72;
parameter character_lowercase_s= 8'h73;
parameter character_lowercase_t= 8'h74;
parameter character_lowercase_u= 8'h75;
parameter character_lowercase_v= 8'h76;
parameter character_lowercase_w= 8'h77;
parameter character_lowercase_x= 8'h78;
parameter character_lowercase_y= 8'h79;
parameter character_lowercase_z= 8'h7A;

//Other Characters
parameter character_colon = 8'h3A;          //':'
parameter character_stop = 8'h2E;           //'.'
parameter character_semi_colon = 8'h3B;   //';'
parameter character_minus = 8'h2D;         //'-'
parameter character_divide = 8'h2F;         //'/'
parameter character_plus = 8'h2B;          //'+'
parameter character_comma = 8'h2C;          // ','
parameter character_less_than = 8'h3C;    //'<'
parameter character_greater_than = 8'h3E; //'>'
parameter character_equals = 8'h3D;         //'='
parameter character_question = 8'h3F;      //'?'
parameter character_dollar = 8'h24;         //'$'
parameter character_space=8'h20;           //' '     
parameter character_exclaim=8'h21;          //'!'


wire Clock_1KHz, Clock_1Hz;
wire Sample_Clk_Signal;

//=======================================================================================================================
//
// Insert your code for Lab2 here!
//
//
wire CLK_22, CLK_22_SYNC; 
wire [31:0] speedometer; //CLOCK wire

wire [7:0] audio_signal;  
//Audio Generation Signal
//Note that the audio needs signed data - so convert 1 bit to 8 bits signed
wire [7:0] audio_data = audio_signal; // = {~Sample_Clk_Signal,{7{Sample_Clk_Signal}}}; //generate signed sample audio signal

wire start, finish;                   // between FSM and ADDRESS_CNTRL
wire play, dir, rst, finish_keyboard; // keyboard wires


wire            flash_mem_read;
wire            flash_mem_waitrequest;
wire    [22:0]  flash_mem_address;
wire    [31:0]  flash_mem_readdata;
wire            flash_mem_readdatavalid;
wire    [3:0]   flash_mem_byteenable = 4'b1111;


COUNTER                           SPEED_CONTROL (.clk(CLK_50M), .up(speed_up_event), .down(speed_down_event), .rst(speed_reset_event),.count(speedometer)); 
//increment, decrement or reset a certain value 
LAB1V2                            CLOCK_DIVIDER (.rst(0), .clk(CLK_50M), .constant(speedometer), .clk_div(CLK_22)); 
//divides clocks based on the given value 
async_trap_and_reset_gen_1_pulse  CLK_22_synchronizer(.async_sig(CLK_22), .outclk(CLK_50M), .out_sync_sig(CLK_22_SYNC), .auto_reset(1'b1), .reset(1'b1));
//synchronizes the 22KHz clock signal
FSM_MEM                           memory_talk1(.clk(CLK_50M), .read(flash_mem_read), .waitrequest(flash_mem_waitrequest), 
                                  .data_valid(flash_mem_readdatavalid), .in(start), .out(finish)); 

ADDRESS_CNTRL                     addr_and_data_manager(.clk(CLK_50M), .frequency_clk(CLK_22_SYNC), 
                                  .play(play), .dir(dir), .rst(rst), //keyboard input signals
                                  .flash_stop(finish), .flash_data(flash_mem_readdata), .flash_begin(start), 
                                  .address(flash_mem_address), .read(flash_mem_read), .finish_keyboard(finish_keyboard),
                                  .out_data(audio_signal)); 
//handles the audio part 
KEYBOARD                          keyboard_cntrl(.clk(CLK_50M), .key(kbd_received_ascii_code), .finish_read(finish_keyboard), .ready(kbd_data_ready), .play(play), .dir(dir), .rst(rst));
//handles keyboard signals 
flash flash_inst (
    .clk_clk                 (CLK_50M),
    .reset_reset_n           (1'b1),
    .flash_mem_write         (1'b0),
    .flash_mem_burstcount    (1'b1),
    .flash_mem_byteenable    (flash_mem_byteenable), //important in
    .flash_mem_read          (flash_mem_read), //important in
    .flash_mem_address       (flash_mem_address), //important in
    .flash_mem_writedata     (), // maybe empty?
    .flash_mem_readdata      (flash_mem_readdata), //important out
    .flash_mem_readdatavalid (flash_mem_readdatavalid), //important out 
    .flash_mem_waitrequest   (flash_mem_waitrequest)// important out 
);
            

assign Sample_Clk_Signal = Clock_1KHz;




//======================================================================================
// 
// Keyboard Interface
//
//

wire ps2c, ps2d; //filtered kbd wires
wire kbd_data_ready, Kbd_to_LCD_finish;

doublesync ps2c_doublsync
(.indata(PS2_CLK),
.outdata(ps2c),
.clk(CLK_50M),
.reset(1'b1));

doublesync ps2d_doublsync
(.indata(PS2_DAT),
.outdata(ps2d),
.clk(CLK_50M),
.reset(1'b1));

wire reset_kbd_data;
(* KEEP = "TRUE" *) wire conv_now_ignore_timing;
 
wire [7:0] kbd_received_ascii_code, kbd_scan_code;
    
Kbd_ctrl Kbd_Controller(
.kbd_clk(ps2c), 
.kbd_data(ps2d),
 .clk(CLK_50M), 
.scan_code(kbd_scan_code), 
.reset_kbd_reg(~reset_kbd_data), 
.data_ready(kbd_data_ready)
);
                
key2ascii kbd2ascii(
.key_code(kbd_scan_code),
.ascii_code(kbd_received_ascii_code),
.clk(conv_now_ignore_timing)
); 
            
parameter scope_info_bytes = 16;
parameter scope_info_bits_per_byte = 8;

wire [15:0] write_kbd_debug;

wire  [scope_info_bits_per_byte-1:0] scope_info0, scope_info1, scope_info2,
     scope_info3, scope_info4, scope_info5, scope_info6, scope_info7, scope_info8, 
     scope_info9, scope_info10, scope_info11, scope_info12, scope_info13, 
     scope_info14, scope_info15;
                
Write_Kbd_To_Scope_LCD Write_Kbd_To_LCD1
(.kbd_ascii_data(kbd_received_ascii_code), 
              .kbd_ready(kbd_data_ready), .reset_kbd_data(reset_kbd_data), 
                     .sm_clk(CLK_50M), .reset(1'b1), 
                     .finish(Kbd_to_LCD_finish), 
                     .scope_info0(scope_info0), 
                     .scope_info1(scope_info1),
                     .scope_info2(scope_info2),
                     .scope_info3(scope_info3),
                     .scope_info4(scope_info4),
                     .scope_info5(scope_info5),
                     .scope_info6(scope_info6),
                     .scope_info7(scope_info7),
                     .scope_info8(scope_info8),
                     .scope_info9(scope_info9),
                     .scope_info10(scope_info10),
                     .scope_info11(scope_info11),
                     .scope_info12(scope_info12),
                     .scope_info13(scope_info13),
                     .scope_info14(scope_info14),
                     .scope_info15(scope_info15),
                     .debug(write_kbd_debug),
                     .convert_now(conv_now_ignore_timing)
    );
                
//=====================================================================================
//
// LCD Scope Acquisition Circuitry Wire Definitions                 
//
//=====================================================================================

wire allow_run_LCD_scope;
wire [15:0] scope_channelA, scope_channelB;
(* keep = 1, preserve = 1 *)wire scope_clk;
reg user_scope_enable_trigger;
wire user_scope_enable;
wire user_scope_enable_trigger_path0, user_scope_enable_trigger_path1;
wire scope_enable_source = SW[8];
wire choose_LCD_or_SCOPE = SW[9];


doublesync user_scope_enable_sync1(.indata(scope_enable_source),
                  .outdata(user_scope_enable),
                  .clk(CLK_50M),
                  .reset(1'b1)); 

//Generate the oscilloscope clock
Generate_Arbitrary_Divided_Clk32 
Generate_LCD_scope_Clk(
.inclk(CLK_50M),
.outclk(scope_clk),
.outclk_Not(),
.div_clk_count(scope_sampling_clock_count),
.Reset(1'h1));

//Scope capture channels
//Scope capture channels

(* keep = 1, preserve = 1 *) logic ScopeChannelASignal;
(* keep = 1, preserve = 1 *) logic ScopeChannelBSignal;

assign ScopeChannelASignal = Sample_Clk_Signal;
assign ScopeChannelBSignal = SW[1];
//Scope capture channels

scope_capture LCD_scope_channelA(
.clk(scope_clk),
.the_signal(ScopeChannelASignal),
.capture_enable(allow_run_LCD_scope & user_scope_enable), 
.captured_data(scope_channelA), //Insert your channel B signal here
.reset(1'b1));

scope_capture LCD_scope_channelB
(
.clk(scope_clk),
.the_signal(ScopeChannelBSignal),
.capture_enable(allow_run_LCD_scope & user_scope_enable), 
.captured_data(scope_channelB), //Insert your channel A signal here
.reset(1'b1));

//The LCD scope and display
LCD_Scope_Encapsulated_pacoblaze_wrapper LCD_LED_scope(
					    //LCD control signals
					    .lcd_d(GPIO_0[7:0]),
					    .lcd_rs(GPIO_0[8]),
					    .lcd_rw(GPIO_0[9]),
					    .lcd_e(GPIO_0[10]),
					    .clk(CLK_50M),
                
                        //LCD Display values
                      .InH(audio_signal),
                      .InG(8'h00),
                      .InF(8'h00),
                      .InE(8'h00),
                      .InD(8'h00),
                      .InC(8'h00),
                      .InB(8'h00),
                      .InA(audio_signal),
                          
                     //LCD display information signals
                         .InfoH({scope_info15,scope_info14}),
                          .InfoG({scope_info13,scope_info12}),
                          .InfoF({scope_info11,scope_info10}),
                          .InfoE({scope_info9,scope_info8}),
                          .InfoD({scope_info7,scope_info6}),
                          .InfoC({scope_info5,scope_info4}),
                          .InfoB({scope_info3,scope_info2}),
                          .InfoA({scope_info1,scope_info0}),
                          
                  //choose to display the values or the oscilloscope
                          .choose_scope_or_LCD(choose_LCD_or_SCOPE),
                          
                  //scope channel declarations
                          .scope_channelA(scope_channelA), //don't touch
                          .scope_channelB(scope_channelB), //don't touch
                          
                  //scope information generation
                          .ScopeInfoA({character_1,character_K,character_H,character_lowercase_z}),
                          .ScopeInfoB({character_S,character_W,character_1,character_space}),
                          
                 //enable_scope is used to freeze the scope just before capturing 
                 //the waveform for display (otherwise the sampling would be unreliable)
                          .enable_scope(allow_run_LCD_scope) //don't touch
                          
    );  
    

//=====================================================================================
//
//  Seven-Segment and speed control
//
//=====================================================================================

wire speed_up_event, speed_down_event;

//Generate 1 KHz Clock
Generate_Arbitrary_Divided_Clk32 
Gen_1KHz_clk
(
.inclk(CLK_50M),
.outclk(Clock_1KHz),
.outclk_Not(),
.div_clk_count(32'h61A6), //change this if necessary to suit your module
.Reset(1'h1)); 

wire speed_up_raw;
wire speed_down_raw;

doublesync 
key0_doublsync
(.indata(!KEY[0]),
.outdata(speed_up_raw),
.clk(Clock_1KHz),
.reset(1'b1));


doublesync 
key1_doublsync
(.indata(!KEY[1]),
.outdata(speed_down_raw),
.clk(Clock_1KHz),
.reset(1'b1));


parameter num_updown_events_per_sec = 10;
parameter num_1KHZ_clocks_between_updown_events = 1000/num_updown_events_per_sec;

reg [15:0] updown_counter = 0;
always @(posedge Clock_1KHz)
begin
      if (updown_counter >= num_1KHZ_clocks_between_updown_events)
      begin
            if (speed_up_raw)
            begin
                  speed_up_event_trigger <= 1;          
            end 
            
            if (speed_down_raw)
            begin
                  speed_down_event_trigger <= 1;            
            end 
            updown_counter <= 0;
      end
      else 
      begin
           updown_counter <= updown_counter + 1;
           speed_up_event_trigger <=0;
           speed_down_event_trigger <= 0;
      end     
end

wire speed_up_event_trigger;
wire speed_down_event_trigger;

async_trap_and_reset_gen_1_pulse 
make_speedup_pulse
(
 .async_sig(speed_up_event_trigger), 
 .outclk(CLK_50M), 
 .out_sync_sig(speed_up_event), 
 .auto_reset(1'b1), 
 .reset(1'b1)
 );
 
async_trap_and_reset_gen_1_pulse 
make_speedown_pulse
(
 .async_sig(speed_down_event_trigger), 
 .outclk(CLK_50M), 
 .out_sync_sig(speed_down_event), 
 .auto_reset(1'b1), 
 .reset(1'b1)
 );


wire speed_reset_event; 

doublesync 
key2_doublsync
(.indata(!KEY[2]),
.outdata(speed_reset_event),
.clk(CLK_50M),
.reset(1'b1));

parameter oscilloscope_speed_step = 100;

wire [15:0] speed_control_val;                      
speed_reg_control 
speed_reg_control_inst
(
.clk(CLK_50M),
.up_event(speed_up_event),
.down_event(speed_down_event),
.reset_event(speed_reset_event),
.speed_control_val(speed_control_val)
);

logic [15:0] scope_sampling_clock_count;
parameter [15:0] default_scope_sampling_clock_count = 12499; //2KHz


always @ (posedge CLK_50M) 
begin
    scope_sampling_clock_count <= default_scope_sampling_clock_count+{{16{speed_control_val[15]}},speed_control_val};
end 

        
        
logic [7:0] Seven_Seg_Val[5:0];
logic [3:0] Seven_Seg_Data[5:0];
    
SevenSegmentDisplayDecoder SevenSegmentDisplayDecoder_inst0(.ssOut(Seven_Seg_Val[0]), .nIn(Seven_Seg_Data[0]));
SevenSegmentDisplayDecoder SevenSegmentDisplayDecoder_inst1(.ssOut(Seven_Seg_Val[1]), .nIn(Seven_Seg_Data[1]));
SevenSegmentDisplayDecoder SevenSegmentDisplayDecoder_inst2(.ssOut(Seven_Seg_Val[2]), .nIn(Seven_Seg_Data[2]));
SevenSegmentDisplayDecoder SevenSegmentDisplayDecoder_inst3(.ssOut(Seven_Seg_Val[3]), .nIn(Seven_Seg_Data[3]));
SevenSegmentDisplayDecoder SevenSegmentDisplayDecoder_inst4(.ssOut(Seven_Seg_Val[4]), .nIn(Seven_Seg_Data[4]));
SevenSegmentDisplayDecoder SevenSegmentDisplayDecoder_inst5(.ssOut(Seven_Seg_Val[5]), .nIn(Seven_Seg_Data[5]));

assign HEX0 = Seven_Seg_Val[0];
assign HEX1 = Seven_Seg_Val[1];
assign HEX2 = Seven_Seg_Val[2];
assign HEX3 = Seven_Seg_Val[3];
assign HEX4 = Seven_Seg_Val[4];
assign HEX5 = Seven_Seg_Val[5];
            
wire Clock_2Hz;
            
Generate_Arbitrary_Divided_Clk32 
Gen_2Hz_clk
(.inclk(CLK_50M),
.outclk(Clock_2Hz),
.outclk_Not(),
.div_clk_count(32'h17D7840 >> 1),
.Reset(1'h1)
); 
        
logic [23:0] actual_7seg_output;
reg [23:0] regd_actual_7seg_output;

always @(posedge Clock_2Hz)
begin
    regd_actual_7seg_output <= actual_7seg_output;
    Clock_1Hz <= ~Clock_1Hz;
end


assign Seven_Seg_Data[0] = regd_actual_7seg_output[3:0];
assign Seven_Seg_Data[1] = regd_actual_7seg_output[7:4];
assign Seven_Seg_Data[2] = regd_actual_7seg_output[11:8];
assign Seven_Seg_Data[3] = regd_actual_7seg_output[15:12];
assign Seven_Seg_Data[4] = regd_actual_7seg_output[19:16];
assign Seven_Seg_Data[5] = regd_actual_7seg_output[23:20];
    
assign actual_7seg_output =  scope_sampling_clock_count;




//=======================================================================================================================
//
//   Audio controller code - do not touch
//
//========================================================================================================================
wire [$size(audio_data)-1:0] actual_audio_data_left, actual_audio_data_right;
wire audio_left_clock, audio_right_clock;

to_slow_clk_interface 
interface_actual_audio_data_right
 (.indata(audio_data),
  .outdata(actual_audio_data_right),
  .inclk(CLK_50M),
  .outclk(audio_right_clock));
   
   
to_slow_clk_interface 
interface_actual_audio_data_left
 (.indata(audio_data),
  .outdata(actual_audio_data_left),
  .inclk(CLK_50M),
  .outclk(audio_left_clock));
   

audio_controller 
audio_control(
  // Clock Input (50 MHz)
  .iCLK_50(CLK_50M), // 50 MHz
  .iCLK_28(), // 27 MHz
  //  7-SEG Displays
  // I2C
  .I2C_SDAT(FPGA_I2C_SDAT), // I2C Data
  .oI2C_SCLK(FPGA_I2C_SCLK), // I2C Clock
  // Audio CODEC
  .AUD_ADCLRCK(AUD_ADCLRCK),                    //  Audio CODEC ADC LR Clock
  .iAUD_ADCDAT(AUD_ADCDAT),                 //  Audio CODEC ADC Data
  .AUD_DACLRCK(AUD_DACLRCK),                    //  Audio CODEC DAC LR Clock
  .oAUD_DACDAT(AUD_DACDAT),                 //  Audio CODEC DAC Data
  .AUD_BCLK(AUD_BCLK),                      //  Audio CODEC Bit-Stream Clock
  .oAUD_XCK(AUD_XCK),                       //  Audio CODEC Chip Clock
  .audio_outL({actual_audio_data_left,8'b1}), 
  .audio_outR({actual_audio_data_right,8'b1}),
  .audio_right_clock(audio_right_clock), 
  .audio_left_clock(audio_left_clock)
);

endmodule
//=======================================================================================================================
//
//   End Audio controller code
//
//========================================================================================================================            
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/*
module sync_machine(in,clk,rst,out); //Syncing for clock input into FSM 
parameter n = 1;
input [n-1:0] in; 
input clk, rst; 
output reg [n-1:0] out; 
reg first, second; 

always@(posedge clk or negedge rst)
    begin 
        if (rst == 1'b0) begin first <= 1'b0; second <= 1'b0; end 
        else             begin first <= in; second <= first; end 
    end 
assign out = second; 
endmodule
////////////////////////////////////////////////////////////////////////////////////////////////
module counterses(clk,limit,rst,count); //Address counter 
parameter n = 32;
input [n-1:0] limit;  
input clk,rst; 
output reg [n-1:0] count; 
reg [n-1:0] counterino; 
always@(posedge clk) 
    begin 
        if(rst)                          begin counterino <= 0; end 
        else if ((counterino != limit) ) begin counterino <= count+1: end
        else if ((counterino == limit) ) begin counterino <= 0; end 
        else                             begin counterino <= counterino; end
    end
assign count = counterino; 
endmodule
/////////////////////////////////////////////////////////////////////////////////////////////// 
module COUNTER(clk, up, down, rst,count); 
 
input up, down, rst, clk; 
output reg [31:0] count; 
 
reg [5:0] state ; 

parameter idle1       = 6'b000000;
parameter idle2       = 6'b000001;
parameter idle3       = 6'b000010;
parameter begin_state = 6'b000100;
parameter up_state    = 6'b001000;
parameter down_state  = 6'b010000;
parameter reset_state = 6'b100000;


always_ff@(posedge clk)
    begin
	    case(state) 
        begin_state:                    state <= idle1; 
	    idle1: 	                        state <= (up)?           up_state   : idle2;
	    idle2:                          state <= (down)?         down_state : idle3; 
        idle3:                          state <= (rst)?          reset_state: idle1;
	    up_state:                       state <=                 idle; 
	    down_state:                     state <=                 idle; 
	    reset_state:                    state <=                 idle; 
	    default:                        state <=                 idle; 
	endcase 
    end
always_ff@(posedge clk)
    begin
	    case(state) 
        begin_state:                    count <= 32'd1136; 
        reset_state:                    count <= 32'd1136; 
	    up_state:                       count <= count + 32'd50; 
	    down_state:                     count <= count - 32'd50; 
	    default:                        count <= count; 
	endcase 
    end

endmodule
*/

module LAB1V2(rst, clk, constant, clk_div); //clock divider code from LAB 1
parameter n= 32;
input clk;  
input rst;
input [n-1:0] constant; 
output reg clk_div = 0; 
reg [n-1:0] counterboy; 
	
always@(posedge clk) 
    begin 
	    if (rst == 1) begin counterboy <= 0; clk_div <= 0; end 
	    else          begin if (counterboy < constant -1) begin counterboy <= counterboy + 1; end 
                            else                          begin counterboy <= 0; clk_div <= ~clk_div; end end 
	end 
endmodule 


module COUNTER(clk, up, down, rst,count); 
 
input up, down, rst, clk; 
output reg [31:0] count; 
reg [31:0 ] counterino = 32'd1136; 
always_ff @(posedge clk)
    begin
        if (rst)    begin counterino <= 32'd1136; end                 //if rst count = 1136
        else if (up) begin counterino <= counterino + 32'd15; end     //if up then count > 1136
        else if (down) begin counterino <= counterino - 32'd15; end   //if down then count < 1136
        else begin counterino <= counterino; end
    end 
assign count = counterino; 
endmodule


module FSM_MEM(clk, read, waitrequest, data_valid, in, out); 
input clk;                                //Trivial
input read, data_valid, waitrequest;      //FROM MEMORY BLOCK 
input in;                              //from ADDRESS_CNTRL
output reg out;                        //to ADDRESS_CNTRL
reg [4:0] state;   //logic [5:0] state; 

parameter idle                         = 5'b0000_0; 
parameter check_oper                   = 5'b0001_0; 
parameter wait_for_waitrequest_negedge = 5'b0010_0; 
parameter wait_for_datavalid_negedge   = 5'b0100_0; 
parameter again                        = 5'b1000_1; 

always_ff@(posedge clk)
    begin
	    case(state) 
	    idle: 	                        state <= (in)?           check_oper : idle;
	    check_oper:                     state <= (read)?         wait_for_waitrequest_negedge : check_oper; 
	    wait_for_waitrequest_negedge:   state <= (~waitrequest)? wait_for_datavalid_negedge : wait_for_datavalid_negedge; 
	    wait_for_datavalid_negedge:     state <= (~data_valid)?  again : wait_for_datavalid_negedge; 
	    again:                          state <=                 idle;
	    default:                        state <=                 idle; 
	endcase 
    end
assign out = state[0]; 
endmodule 


module ADDRESS_CNTRL(clk, frequency_clk, play, dir, rst, flash_stop, flash_data, flash_begin, address, read, finish_keyboard, out_data); 

input clk, frequency_clk;  //trivial
input play, dir, rst;      //from Keyboard
input flash_stop;          //from FSM_MEM
input [31:0] flash_data;   //from flash memory 

output flash_begin, finish_keyboard, read; // to FSM_MEM // to KEYBOARD // to falsh memory 
output [22:0] address; //to flash memory 
output [7:0] out_data; //To audio 
reg [10:0] state;   //logic [5:0] state;

parameter idle_state                = 11'b000000000_00; 
parameter read_state                = 11'b000000001_01; 
parameter wait_to_read_lower_bits   = 11'b000000010_00; 
parameter read_lower_bits           = 11'b000000100_00; 
parameter wait_to_read_upper_bits   = 11'b000001000_00; 
parameter read_upper_bits           = 11'b000010000_00; 
parameter check_oper_keyboard       = 11'b000100000_00; 
parameter minus_speed               = 11'b001000000_00; 
parameter plus_speed                = 11'b010000000_00; 
parameter again                     = 11'b100000000_10; 


///////SEQUENTIAL
always_ff@(posedge clk) 
    begin 
	    case(state) 
		idle_state:                 state <= ((play)?            read_state : idle_state); 
		read_state:                 state <= ((flash_stop)?      wait_to_read_lower_bits: read_state);   
		wait_to_read_lower_bits:    state <= ((frequency_clk)?   read_lower_bits : wait_to_read_lower_bits); 
		read_lower_bits:            state <=                     wait_to_read_upper_bits; 
		wait_to_read_upper_bits:    state <= ((frequency_clk)?   read_upper_bits : wait_to_read_upper_bits);   
		read_upper_bits:            state <=                     check_oper_keyboard;
        check_oper_keyboard:        state <= ((dir)?             minus_speed : plus_speed);
		plus_speed:                 state <= again; 
		minus_speed:                state <= again;  
		again:                      state <= idle_state; 
		default:                    state <= idle_state; 	
	    endcase 
    end 
///////OUTPUTS
    assign flash_begin = state[0]; 
    assign read = state[0]; 
    assign finish_keyboard = state[1]; 

always_ff@(posedge clk) 
    begin 
	    case (state)
	    read_lower_bits:begin out_data <= ((dir)? flash_data[31:24]: flash_data[15:8] ); address <= address; end
        read_upper_bits:begin out_data <= ((dir)? flash_data[15:8] : flash_data[31:24]); address <= address; end
        minus_speed:
                    begin 
                    if(rst) begin address <= 23'h7FFFF;out_data <= out_data; end	    
			        else if (address == 0) begin address <= 23'h7FFFF;out_data <= out_data;end
			        else begin address <= address - 23'd1;out_data <= out_data;end 	
			        end 	
	    plus_speed:
                    begin  
			        if(rst) begin address <= 0;out_data <= out_data; end	    
			        else if (address == 23'h7FFFF) begin address <= 0;out_data <= out_data;end
			        else begin address <= address + 23'd1;out_data <= out_data;end 	  
			        end 
	    default: begin address <= address; out_data <= out_data; end
	    endcase 
    end 

endmodule 



module KEYBOARD(clk,  ready, finish_read, key, play, dir, rst);
input clk, finish_read, ready;
input [7:0] key; 
output play, rst, dir; 
reg [8:0] state; 

parameter check_keyboard = 9'b000000_000; //play/rst/dir
parameter normal_rst     = 9'b000010_110;
parameter normal         = 9'b000001_100;
parameter normal_pause   = 9'b000100_000;
parameter backward_rst   = 9'b010000_111;
parameter backward       = 9'b001000_101;
parameter backward_pause = 9'b100000_000;

//Uppercase Letters

parameter character_B =8'h42;
parameter character_D =8'h44;
parameter character_E =8'h45;
parameter character_F =8'h46;
parameter character_R =8'h52;


assign play = state[2]; 
assign rst = state[1]; 
assign dir = state[0]; 

	
	
always_ff@(posedge clk)
    begin
		case(state)
        normal_rst: 					      state <= finish_read? normal: normal_rst;
        backward_rst: 					      state <= finish_read? backward: backward_rst;
		check_keyboard: 
            begin 
			if      (key == character_E) state <= normal; 
            else if (key == character_F) state <= normal_pause;
			else if (key == character_B) state <= backward_pause; 
			else                         state <= check_keyboard; 
			end 
		normal: 
            begin 
			if     (key == character_R) begin state <= ready? normal_rst : normal; end 
            else if(key == character_B) begin state <= backward; end 
			else if(key == character_D) begin state <= normal_pause; end
			else                              state <= normal; 
			end 	
		normal_pause:
            begin 
			if      (key == character_R) begin state <= normal_rst; end 
            else if (key == character_B) begin state <= backward_pause; end
			else if (key == character_E) begin state <= normal; end
	        else                               state <= normal_pause; 
			end 
		backward: 
            begin 
			if     (key == character_R) begin state <= ready? backward_rst : backward; end 
            else if(key == character_F) begin state <= normal; end 
			else if(key == character_D) begin state <= backward_pause; end
			else                              state <= backward; 
			end 	
		backward_pause:
            begin 
			if      (key == character_R) begin state <= backward_rst; end 
			else if (key == character_F) begin state <= normal_pause; end
			else if (key == character_E) begin state <= backward; end
	        else                               state <= backward_pause; 
			end 
		default: state <= check_keyboard; 
		endcase
	end
endmodule


